-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.0 Build 156 04/24/2013 SJ Web Edition
-- Created on Tue Apr 30 20:03:37 2019

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY moor IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        N : IN STD_LOGIC := '0';
        D : IN STD_LOGIC := '0';
        R : OUT STD_LOGIC
    );
END moor;

ARCHITECTURE BEHAVIOR OF moor IS
    TYPE type_fstate IS (S0,S1,S2,S3,S4);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,N,D)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= S0;
            R <= '0';
        ELSE
            R <= '0';
            CASE fstate IS
                WHEN S0 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= S1;
                    ELSIF (((D = '1') AND NOT((N = '1')))) THEN
                        reg_fstate <= S0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S0;
                    END IF;
                WHEN S1 =>
                    IF ((D = '1')) THEN
                        reg_fstate <= S2;
                    ELSIF (((N = '1') AND NOT((D = '1')))) THEN
                        reg_fstate <= S1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S1;
                    END IF;
                WHEN S2 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= S3;
                    ELSIF (((D = '1') AND NOT((N = '1')))) THEN
                        reg_fstate <= S0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S2;
                    END IF;
                WHEN S3 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= S4;
                    ELSIF (((D = '1') AND NOT((N = '1')))) THEN
                        reg_fstate <= S0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= S3;
                    END IF;
                WHEN S4 =>
                    reg_fstate <= S0;

                    R <= '1';
                WHEN OTHERS => 
                    R <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
