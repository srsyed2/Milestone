// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.0 Build 156 04/24/2013 SJ Web Edition
// Created on Tue Apr 30 19:57:51 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module moor (
    clock,reset,N,D,
    R);

    input clock;
    input reset;
    input N;
    input D;
    tri0 reset;
    tri0 N;
    tri0 D;
    output R;
    reg R;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter S0=0,S1=1,S2=2,S3=3,S4=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or N or D)
    begin
        if (reset) begin
            reg_fstate <= S0;
            R <= 1'b0;
        end
        else begin
            R <= 1'b0;
            case (fstate)
                S0: begin
                    if (N)
                        reg_fstate <= S1;
                    else if ((D & ~(N)))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S0;
                end
                S1: begin
                    if (D)
                        reg_fstate <= S2;
                    else if ((N & ~(D)))
                        reg_fstate <= S1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S1;
                end
                S2: begin
                    if (N)
                        reg_fstate <= S3;
                    else if ((D & ~(N)))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S2;
                end
                S3: begin
                    if (N)
                        reg_fstate <= S4;
                    else if ((D & ~(N)))
                        reg_fstate <= S0;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= S3;
                end
                S4: begin
                    reg_fstate <= S0;

                    R <= 1'b1;
                end
                default: begin
                    R <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // moor
