// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 13.0.0 Build 156 04/24/2013 SJ Web Edition
// Created on Sun Apr 21 17:55:47 2019

// synthesis message_off 10175

`timescale 1ns/1ns

module vendingmoore (
    reset,clock,N,D,
    R);

    input reset;
    input clock;
    input N;
    input D;
    tri0 reset;
    tri0 N;
    tri0 D;
    output R;
    reg R;
    reg [4:0] fstate;
    reg [4:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or N or D)
    begin
        if (reset) begin
            reg_fstate <= state1;
            R <= 1'b0;
        end
        else begin
            R <= 1'b0;
            case (fstate)
                state1: begin
                    if (N)
                        reg_fstate <= state2;
                    else if ((D & ~(N)))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    if (D)
                        reg_fstate <= state3;
                    else if ((N & ~(D)))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;
                end
                state3: begin
                    if (N)
                        reg_fstate <= state4;
                    else if ((D & ~(N)))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;
                end
                state4: begin
                    if (N)
                        reg_fstate <= state5;
                    else if ((D & ~(N)))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;
                end
                state5: begin
                    reg_fstate <= state1;

                    R <= 1'b1;
                end
                default: begin
                    R <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // vendingmoore
